package pack2;
import pack1 :: pp1;
import pack1 :: pp2;
export pack1:: *;
export pack1:: *;
endpackage