package pack1;

parameter       pp1 = 10 ;
parameter       pp2 = 20 ;
integer         i   ;
byte            b   ;
endpackage