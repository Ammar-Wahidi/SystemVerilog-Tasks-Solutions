`define M1(a,b) \
initial \
        begin \
            $display(a); \
            $display(b); \
        end 

`define M2 30 
`define plus(a,b) a+b
