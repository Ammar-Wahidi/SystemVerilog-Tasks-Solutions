package Memory_package_UVM;

import uvm_pkg::*;
`include "uvm_macros.svh"
`include "my_sequence_item.svh"
`include "my_sequence.svh"
`include "my_sequence_rand.svh"
`include "my_sequencer.svh"
`include "my_driver.svh"
`include "my_monitor.svh"
`include "my_subscriber.svh"
`include "my_scoreboard.svh"
`include "my_agent.svh"
`include "my_env.svh"
`include "my_test.svh"

endpackage