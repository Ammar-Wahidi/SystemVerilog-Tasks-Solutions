module top();
import uvm_pkg ::* ;
import pack1 ::* ;

initial
begin
    run_test("my_test") ;
end  
endmodule