package pack3;
import pack2::*;
export pack2:: pp1;
export pack2:: pp2;
endpackage